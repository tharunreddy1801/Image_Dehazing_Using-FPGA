module ADD(
input [15:0]a,
input [31:0]b,
output [31:0]sum
);
assign sum = a + b;
endmodule