module ATM_LUT (
    input  [7:0] in_val,
    output reg [15:0] out_val
);

always @(*) begin
    case (in_val)
        8'd  1: out_val = 16'd65535;  // 1/1 ? 1.00000000
        8'd  2: out_val = 16'd32768;  // 1/2 ? 0.50000000
        8'd  3: out_val = 16'd21845;  // 1/3 ? 0.33333333
        8'd  4: out_val = 16'd16384;  // 1/4 ? 0.25000000
        8'd  5: out_val = 16'd13107;  // 1/5 ? 0.20000000
        8'd  6: out_val = 16'd10923;  // 1/6 ? 0.16666667
        8'd  7: out_val = 16'd 9362;  // 1/7 ? 0.14285714
        8'd  8: out_val = 16'd 8192;  // 1/8 ? 0.12500000
        8'd  9: out_val = 16'd 7282;  // 1/9 ? 0.11111111
        8'd 10: out_val = 16'd 6554;  // 1/10 ? 0.10000000
        8'd 11: out_val = 16'd 5958;  // 1/11 ? 0.09090909
        8'd 12: out_val = 16'd 5461;  // 1/12 ? 0.08333333
        8'd 13: out_val = 16'd 5041;  // 1/13 ? 0.07692308
        8'd 14: out_val = 16'd 4681;  // 1/14 ? 0.07142857
        8'd 15: out_val = 16'd 4369;  // 1/15 ? 0.06666667
        8'd 16: out_val = 16'd 4096;  // 1/16 ? 0.06250000
        8'd 17: out_val = 16'd 3855;  // 1/17 ? 0.05882353
        8'd 18: out_val = 16'd 3641;  // 1/18 ? 0.05555556
        8'd 19: out_val = 16'd 3449;  // 1/19 ? 0.05263158
        8'd 20: out_val = 16'd 3277;  // 1/20 ? 0.05000000
        8'd 21: out_val = 16'd 3121;  // 1/21 ? 0.04761905
        8'd 22: out_val = 16'd 2979;  // 1/22 ? 0.04545455
        8'd 23: out_val = 16'd 2849;  // 1/23 ? 0.04347826
        8'd 24: out_val = 16'd 2731;  // 1/24 ? 0.04166667
        8'd 25: out_val = 16'd 2621;  // 1/25 ? 0.04000000
        8'd 26: out_val = 16'd 2521;  // 1/26 ? 0.03846154
        8'd 27: out_val = 16'd 2427;  // 1/27 ? 0.03703704
        8'd 28: out_val = 16'd 2341;  // 1/28 ? 0.03571429
        8'd 29: out_val = 16'd 2260;  // 1/29 ? 0.03448276
        8'd 30: out_val = 16'd 2185;  // 1/30 ? 0.03333333
        8'd 31: out_val = 16'd 2114;  // 1/31 ? 0.03225806
        8'd 32: out_val = 16'd 2048;  // 1/32 ? 0.03125000
        8'd 33: out_val = 16'd 1986;  // 1/33 ? 0.03030303
        8'd 34: out_val = 16'd 1928;  // 1/34 ? 0.02941176
        8'd 35: out_val = 16'd 1872;  // 1/35 ? 0.02857143
        8'd 36: out_val = 16'd 1820;  // 1/36 ? 0.02777778
        8'd 37: out_val = 16'd 1771;  // 1/37 ? 0.02702703
        8'd 38: out_val = 16'd 1725;  // 1/38 ? 0.02631579
        8'd 39: out_val = 16'd 1680;  // 1/39 ? 0.02564103
        8'd 40: out_val = 16'd 1638;  // 1/40 ? 0.02500000
        8'd 41: out_val = 16'd 1598;  // 1/41 ? 0.02439024
        8'd 42: out_val = 16'd 1560;  // 1/42 ? 0.02380952
        8'd 43: out_val = 16'd 1524;  // 1/43 ? 0.02325581
        8'd 44: out_val = 16'd 1489;  // 1/44 ? 0.02272727
        8'd 45: out_val = 16'd 1456;  // 1/45 ? 0.02222222
        8'd 46: out_val = 16'd 1425;  // 1/46 ? 0.02173913
        8'd 47: out_val = 16'd 1394;  // 1/47 ? 0.02127660
        8'd 48: out_val = 16'd 1365;  // 1/48 ? 0.02083333
        8'd 49: out_val = 16'd 1337;  // 1/49 ? 0.02040816
        8'd 50: out_val = 16'd 1311;  // 1/50 ? 0.02000000
        8'd 51: out_val = 16'd 1285;  // 1/51 ? 0.01960784
        8'd 52: out_val = 16'd 1260;  // 1/52 ? 0.01923077
        8'd 53: out_val = 16'd 1237;  // 1/53 ? 0.01886792
        8'd 54: out_val = 16'd 1214;  // 1/54 ? 0.01851852
        8'd 55: out_val = 16'd 1192;  // 1/55 ? 0.01818182
        8'd 56: out_val = 16'd 1170;  // 1/56 ? 0.01785714
        8'd 57: out_val = 16'd 1150;  // 1/57 ? 0.01754386
        8'd 58: out_val = 16'd 1130;  // 1/58 ? 0.01724138
        8'd 59: out_val = 16'd 1111;  // 1/59 ? 0.01694915
        8'd 60: out_val = 16'd 1092;  // 1/60 ? 0.01666667
        8'd 61: out_val = 16'd 1074;  // 1/61 ? 0.01639344
        8'd 62: out_val = 16'd 1057;  // 1/62 ? 0.01612903
        8'd 63: out_val = 16'd 1040;  // 1/63 ? 0.01587302
        8'd 64: out_val = 16'd 1024;  // 1/64 ? 0.01562500
        8'd 65: out_val = 16'd 1008;  // 1/65 ? 0.01538462
        8'd 66: out_val = 16'd  993;  // 1/66 ? 0.01515152
        8'd 67: out_val = 16'd  978;  // 1/67 ? 0.01492537
        8'd 68: out_val = 16'd  964;  // 1/68 ? 0.01470588
        8'd 69: out_val = 16'd  950;  // 1/69 ? 0.01449275
        8'd 70: out_val = 16'd  936;  // 1/70 ? 0.01428571
        8'd 71: out_val = 16'd  923;  // 1/71 ? 0.01408451
        8'd 72: out_val = 16'd  910;  // 1/72 ? 0.01388889
        8'd 73: out_val = 16'd  898;  // 1/73 ? 0.01369863
        8'd 74: out_val = 16'd  886;  // 1/74 ? 0.01351351
        8'd 75: out_val = 16'd  874;  // 1/75 ? 0.01333333
        8'd 76: out_val = 16'd  862;  // 1/76 ? 0.01315789
        8'd 77: out_val = 16'd  851;  // 1/77 ? 0.01298701
        8'd 78: out_val = 16'd  840;  // 1/78 ? 0.01282051
        8'd 79: out_val = 16'd  830;  // 1/79 ? 0.01265823
        8'd 80: out_val = 16'd  819;  // 1/80 ? 0.01250000
        8'd 81: out_val = 16'd  809;  // 1/81 ? 0.01234568
        8'd 82: out_val = 16'd  799;  // 1/82 ? 0.01219512
        8'd 83: out_val = 16'd  790;  // 1/83 ? 0.01204819
        8'd 84: out_val = 16'd  780;  // 1/84 ? 0.01190476
        8'd 85: out_val = 16'd  771;  // 1/85 ? 0.01176471
        8'd 86: out_val = 16'd  762;  // 1/86 ? 0.01162791
        8'd 87: out_val = 16'd  753;  // 1/87 ? 0.01149425
        8'd 88: out_val = 16'd  745;  // 1/88 ? 0.01136364
        8'd 89: out_val = 16'd  736;  // 1/89 ? 0.01123596
        8'd 90: out_val = 16'd  728;  // 1/90 ? 0.01111111
        8'd 91: out_val = 16'd  720;  // 1/91 ? 0.01098901
        8'd 92: out_val = 16'd  712;  // 1/92 ? 0.01086957
        8'd 93: out_val = 16'd  705;  // 1/93 ? 0.01075269
        8'd 94: out_val = 16'd  697;  // 1/94 ? 0.01063830
        8'd 95: out_val = 16'd  690;  // 1/95 ? 0.01052632
        8'd 96: out_val = 16'd  683;  // 1/96 ? 0.01041667
        8'd 97: out_val = 16'd  676;  // 1/97 ? 0.01030928
        8'd 98: out_val = 16'd  669;  // 1/98 ? 0.01020408
        8'd 99: out_val = 16'd  662;  // 1/99 ? 0.01010101
        8'd100: out_val = 16'd  655;  // 1/100 ? 0.01000000
        8'd101: out_val = 16'd  649;  // 1/101 ? 0.00990099
        8'd102: out_val = 16'd  643;  // 1/102 ? 0.00980392
        8'd103: out_val = 16'd  636;  // 1/103 ? 0.00970874
        8'd104: out_val = 16'd  630;  // 1/104 ? 0.00961538
        8'd105: out_val = 16'd  624;  // 1/105 ? 0.00952381
        8'd106: out_val = 16'd  618;  // 1/106 ? 0.00943396
        8'd107: out_val = 16'd  612;  // 1/107 ? 0.00934579
        8'd108: out_val = 16'd  607;  // 1/108 ? 0.00925926
        8'd109: out_val = 16'd  601;  // 1/109 ? 0.00917431
        8'd110: out_val = 16'd  596;  // 1/110 ? 0.00909091
        8'd111: out_val = 16'd  590;  // 1/111 ? 0.00900901
        8'd112: out_val = 16'd  585;  // 1/112 ? 0.00892857
        8'd113: out_val = 16'd  580;  // 1/113 ? 0.00884956
        8'd114: out_val = 16'd  575;  // 1/114 ? 0.00877193
        8'd115: out_val = 16'd  570;  // 1/115 ? 0.00869565
        8'd116: out_val = 16'd  565;  // 1/116 ? 0.00862069
        8'd117: out_val = 16'd  560;  // 1/117 ? 0.00854701
        8'd118: out_val = 16'd  555;  // 1/118 ? 0.00847458
        8'd119: out_val = 16'd  551;  // 1/119 ? 0.00840336
        8'd120: out_val = 16'd  546;  // 1/120 ? 0.00833333
        8'd121: out_val = 16'd  542;  // 1/121 ? 0.00826446
        8'd122: out_val = 16'd  537;  // 1/122 ? 0.00819672
        8'd123: out_val = 16'd  533;  // 1/123 ? 0.00813008
        8'd124: out_val = 16'd  529;  // 1/124 ? 0.00806452
        8'd125: out_val = 16'd  524;  // 1/125 ? 0.00800000
        8'd126: out_val = 16'd  520;  // 1/126 ? 0.00793651
        8'd127: out_val = 16'd  516;  // 1/127 ? 0.00787402
        8'd128: out_val = 16'd  512;  // 1/128 ? 0.00781250
        8'd129: out_val = 16'd  508;  // 1/129 ? 0.00775194
        8'd130: out_val = 16'd  504;  // 1/130 ? 0.00769231
        8'd131: out_val = 16'd  500;  // 1/131 ? 0.00763359
        8'd132: out_val = 16'd  496;  // 1/132 ? 0.00757576
        8'd133: out_val = 16'd  493;  // 1/133 ? 0.00751880
        8'd134: out_val = 16'd  489;  // 1/134 ? 0.00746269
        8'd135: out_val = 16'd  485;  // 1/135 ? 0.00740741
        8'd136: out_val = 16'd  482;  // 1/136 ? 0.00735294
        8'd137: out_val = 16'd  478;  // 1/137 ? 0.00729927
        8'd138: out_val = 16'd  475;  // 1/138 ? 0.00724638
        8'd139: out_val = 16'd  471;  // 1/139 ? 0.00719424
        8'd140: out_val = 16'd  468;  // 1/140 ? 0.00714286
        8'd141: out_val = 16'd  465;  // 1/141 ? 0.00709220
        8'd142: out_val = 16'd  462;  // 1/142 ? 0.00704225
        8'd143: out_val = 16'd  458;  // 1/143 ? 0.00699301
        8'd144: out_val = 16'd  455;  // 1/144 ? 0.00694444
        8'd145: out_val = 16'd  452;  // 1/145 ? 0.00689655
        8'd146: out_val = 16'd  449;  // 1/146 ? 0.00684932
        8'd147: out_val = 16'd  446;  // 1/147 ? 0.00680272
        8'd148: out_val = 16'd  443;  // 1/148 ? 0.00675676
        8'd149: out_val = 16'd  440;  // 1/149 ? 0.00671141
        8'd150: out_val = 16'd  437;  // 1/150 ? 0.00666667
        8'd151: out_val = 16'd  434;  // 1/151 ? 0.00662252
        8'd152: out_val = 16'd  431;  // 1/152 ? 0.00657895
        8'd153: out_val = 16'd  428;  // 1/153 ? 0.00653595
        8'd154: out_val = 16'd  426;  // 1/154 ? 0.00649351
        8'd155: out_val = 16'd  423;  // 1/155 ? 0.00645161
        8'd156: out_val = 16'd  420;  // 1/156 ? 0.00641026
        8'd157: out_val = 16'd  417;  // 1/157 ? 0.00636943
        8'd158: out_val = 16'd  415;  // 1/158 ? 0.00632911
        8'd159: out_val = 16'd  412;  // 1/159 ? 0.00628931
        8'd160: out_val = 16'd  410;  // 1/160 ? 0.00625000
        8'd161: out_val = 16'd  407;  // 1/161 ? 0.00621118
        8'd162: out_val = 16'd  405;  // 1/162 ? 0.00617284
        8'd163: out_val = 16'd  402;  // 1/163 ? 0.00613497
        8'd164: out_val = 16'd  400;  // 1/164 ? 0.00609756
        8'd165: out_val = 16'd  397;  // 1/165 ? 0.00606061
        8'd166: out_val = 16'd  395;  // 1/166 ? 0.00602410
        8'd167: out_val = 16'd  392;  // 1/167 ? 0.00598802
        8'd168: out_val = 16'd  390;  // 1/168 ? 0.00595238
        8'd169: out_val = 16'd  388;  // 1/169 ? 0.00591716
        8'd170: out_val = 16'd  386;  // 1/170 ? 0.00588235
        8'd171: out_val = 16'd  383;  // 1/171 ? 0.00584795
        8'd172: out_val = 16'd  381;  // 1/172 ? 0.00581395
        8'd173: out_val = 16'd  379;  // 1/173 ? 0.00578035
        8'd174: out_val = 16'd  377;  // 1/174 ? 0.00574713
        8'd175: out_val = 16'd  374;  // 1/175 ? 0.00571429
        8'd176: out_val = 16'd  372;  // 1/176 ? 0.00568182
        8'd177: out_val = 16'd  370;  // 1/177 ? 0.00564972
        8'd178: out_val = 16'd  368;  // 1/178 ? 0.00561798
        8'd179: out_val = 16'd  366;  // 1/179 ? 0.00558659
        8'd180: out_val = 16'd  364;  // 1/180 ? 0.00555556
        8'd181: out_val = 16'd  362;  // 1/181 ? 0.00552486
        8'd182: out_val = 16'd  360;  // 1/182 ? 0.00549451
        8'd183: out_val = 16'd  358;  // 1/183 ? 0.00546448
        8'd184: out_val = 16'd  356;  // 1/184 ? 0.00543478
        8'd185: out_val = 16'd  354;  // 1/185 ? 0.00540541
        8'd186: out_val = 16'd  352;  // 1/186 ? 0.00537634
        8'd187: out_val = 16'd  350;  // 1/187 ? 0.00534759
        8'd188: out_val = 16'd  349;  // 1/188 ? 0.00531915
        8'd189: out_val = 16'd  347;  // 1/189 ? 0.00529101
        8'd190: out_val = 16'd  345;  // 1/190 ? 0.00526316
        8'd191: out_val = 16'd  343;  // 1/191 ? 0.00523560
        8'd192: out_val = 16'd  341;  // 1/192 ? 0.00520833
        8'd193: out_val = 16'd  340;  // 1/193 ? 0.00518135
        8'd194: out_val = 16'd  338;  // 1/194 ? 0.00515464
        8'd195: out_val = 16'd  336;  // 1/195 ? 0.00512821
        8'd196: out_val = 16'd  334;  // 1/196 ? 0.00510204
        8'd197: out_val = 16'd  333;  // 1/197 ? 0.00507614
        8'd198: out_val = 16'd  331;  // 1/198 ? 0.00505051
        8'd199: out_val = 16'd  329;  // 1/199 ? 0.00502513
        8'd200: out_val = 16'd  328;  // 1/200 ? 0.00500000
        8'd201: out_val = 16'd  326;  // 1/201 ? 0.00497512
        8'd202: out_val = 16'd  324;  // 1/202 ? 0.00495050
        8'd203: out_val = 16'd  323;  // 1/203 ? 0.00492611
        8'd204: out_val = 16'd  321;  // 1/204 ? 0.00490196
        8'd205: out_val = 16'd  320;  // 1/205 ? 0.00487805
        8'd206: out_val = 16'd  318;  // 1/206 ? 0.00485437
        8'd207: out_val = 16'd  317;  // 1/207 ? 0.00483092
        8'd208: out_val = 16'd  315;  // 1/208 ? 0.00480769
        8'd209: out_val = 16'd  314;  // 1/209 ? 0.00478469
        8'd210: out_val = 16'd  312;  // 1/210 ? 0.00476190
        8'd211: out_val = 16'd  311;  // 1/211 ? 0.00473934
        8'd212: out_val = 16'd  309;  // 1/212 ? 0.00471698
        8'd213: out_val = 16'd  308;  // 1/213 ? 0.00469484
        8'd214: out_val = 16'd  306;  // 1/214 ? 0.00467290
        8'd215: out_val = 16'd  305;  // 1/215 ? 0.00465116
        8'd216: out_val = 16'd  303;  // 1/216 ? 0.00462963
        8'd217: out_val = 16'd  302;  // 1/217 ? 0.00460829
        8'd218: out_val = 16'd  301;  // 1/218 ? 0.00458716
        8'd219: out_val = 16'd  299;  // 1/219 ? 0.00456621
        8'd220: out_val = 16'd  298;  // 1/220 ? 0.00454545
        8'd221: out_val = 16'd  297;  // 1/221 ? 0.00452489
        8'd222: out_val = 16'd  295;  // 1/222 ? 0.00450450
        8'd223: out_val = 16'd  294;  // 1/223 ? 0.00448430
        8'd224: out_val = 16'd  293;  // 1/224 ? 0.00446429
        8'd225: out_val = 16'd  291;  // 1/225 ? 0.00444444
        8'd226: out_val = 16'd  290;  // 1/226 ? 0.00442478
        8'd227: out_val = 16'd  289;  // 1/227 ? 0.00440529
        8'd228: out_val = 16'd  287;  // 1/228 ? 0.00438596
        8'd229: out_val = 16'd  286;  // 1/229 ? 0.00436681
        8'd230: out_val = 16'd  285;  // 1/230 ? 0.00434783
        8'd231: out_val = 16'd  284;  // 1/231 ? 0.00432900
        8'd232: out_val = 16'd  282;  // 1/232 ? 0.00431034
        8'd233: out_val = 16'd  281;  // 1/233 ? 0.00429185
        8'd234: out_val = 16'd  280;  // 1/234 ? 0.00427350
        8'd235: out_val = 16'd  279;  // 1/235 ? 0.00425532
        8'd236: out_val = 16'd  278;  // 1/236 ? 0.00423729
        8'd237: out_val = 16'd  277;  // 1/237 ? 0.00421941
        8'd238: out_val = 16'd  275;  // 1/238 ? 0.00420168
        8'd239: out_val = 16'd  274;  // 1/239 ? 0.00418410
        8'd240: out_val = 16'd  273;  // 1/240 ? 0.00416667
        8'd241: out_val = 16'd  272;  // 1/241 ? 0.00414938
        8'd242: out_val = 16'd  271;  // 1/242 ? 0.00413223
        8'd243: out_val = 16'd  270;  // 1/243 ? 0.00411523
        8'd244: out_val = 16'd  269;  // 1/244 ? 0.00409836
        8'd245: out_val = 16'd  267;  // 1/245 ? 0.00408163
        8'd246: out_val = 16'd  266;  // 1/246 ? 0.00406504
        8'd247: out_val = 16'd  265;  // 1/247 ? 0.00404858
        8'd248: out_val = 16'd  264;  // 1/248 ? 0.00403226
        8'd249: out_val = 16'd  263;  // 1/249 ? 0.00401606
        8'd250: out_val = 16'd  262;  // 1/250 ? 0.00400000
        8'd251: out_val = 16'd  261;  // 1/251 ? 0.00398406
        8'd252: out_val = 16'd  260;  // 1/252 ? 0.00396825
        8'd253: out_val = 16'd  259;  // 1/253 ? 0.00395257
        8'd254: out_val = 16'd  258;  // 1/254 ? 0.00393701
        8'd255: out_val = 16'd  257;  // 1/255 ? 0.00392157
        default: out_val = 16'd0;  // undefined for 0
    endcase
end

endmodule