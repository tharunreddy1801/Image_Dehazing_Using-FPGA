module power_luts(
    input wire [7:0] x,
    input wire [7:0] y,
    output reg [15:0] x_pow_03,
    output reg [15:0] y_pow_07
);

always @(*) begin
    case(x)
        8'd0: x_pow_03 = 16'd0;
        8'd1: x_pow_03 = 16'd49;
        8'd2: x_pow_03 = 16'd60;
        8'd3: x_pow_03 = 16'd68;
        8'd4: x_pow_03 = 16'd74;
        8'd5: x_pow_03 = 16'd79;
        8'd6: x_pow_03 = 16'd83;
        8'd7: x_pow_03 = 16'd87;
        8'd8: x_pow_03 = 16'd91;
        8'd9: x_pow_03 = 16'd94;
        8'd10: x_pow_03 = 16'd97;
        8'd11: x_pow_03 = 16'd100;
        8'd12: x_pow_03 = 16'd102;
        8'd13: x_pow_03 = 16'd105;
        8'd14: x_pow_03 = 16'd107;
        8'd15: x_pow_03 = 16'd109;
        8'd16: x_pow_03 = 16'd112;
        8'd17: x_pow_03 = 16'd114;
        8'd18: x_pow_03 = 16'd116;
        8'd19: x_pow_03 = 16'd117;
        8'd20: x_pow_03 = 16'd119;
        8'd21: x_pow_03 = 16'd121;
        8'd22: x_pow_03 = 16'd123;
        8'd23: x_pow_03 = 16'd124;
        8'd24: x_pow_03 = 16'd126;
        8'd25: x_pow_03 = 16'd128;
        8'd26: x_pow_03 = 16'd129;
        8'd27: x_pow_03 = 16'd131;
        8'd28: x_pow_03 = 16'd132;
        8'd29: x_pow_03 = 16'd133;
        8'd30: x_pow_03 = 16'd135;
        8'd31: x_pow_03 = 16'd136;
        8'd32: x_pow_03 = 16'd137;
        8'd33: x_pow_03 = 16'd139;
        8'd34: x_pow_03 = 16'd140;
        8'd35: x_pow_03 = 16'd141;
        8'd36: x_pow_03 = 16'd142;
        8'd37: x_pow_03 = 16'd143;
        8'd38: x_pow_03 = 16'd145;
        8'd39: x_pow_03 = 16'd146;
        8'd40: x_pow_03 = 16'd147;
        8'd41: x_pow_03 = 16'd148;
        8'd42: x_pow_03 = 16'd149;
        8'd43: x_pow_03 = 16'd150;
        8'd44: x_pow_03 = 16'd151;
        8'd45: x_pow_03 = 16'd152;
        8'd46: x_pow_03 = 16'd153;
        8'd47: x_pow_03 = 16'd154;
        8'd48: x_pow_03 = 16'd155;
        8'd49: x_pow_03 = 16'd156;
        8'd50: x_pow_03 = 16'd157;
        8'd51: x_pow_03 = 16'd158;
        8'd52: x_pow_03 = 16'd159;
        8'd53: x_pow_03 = 16'd160;
        8'd54: x_pow_03 = 16'd161;
        8'd55: x_pow_03 = 16'd162;
        8'd56: x_pow_03 = 16'd162;
        8'd57: x_pow_03 = 16'd163;
        8'd58: x_pow_03 = 16'd164;
        8'd59: x_pow_03 = 16'd165;
        8'd60: x_pow_03 = 16'd166;
        8'd61: x_pow_03 = 16'd167;
        8'd62: x_pow_03 = 16'd167;
        8'd63: x_pow_03 = 16'd168;
        8'd64: x_pow_03 = 16'd169;
        8'd65: x_pow_03 = 16'd170;
        8'd66: x_pow_03 = 16'd171;
        8'd67: x_pow_03 = 16'd171;
        8'd68: x_pow_03 = 16'd172;
        8'd69: x_pow_03 = 16'd173;
        8'd70: x_pow_03 = 16'd174;
        8'd71: x_pow_03 = 16'd174;
        8'd72: x_pow_03 = 16'd175;
        8'd73: x_pow_03 = 16'd176;
        8'd74: x_pow_03 = 16'd177;
        8'd75: x_pow_03 = 16'd177;
        8'd76: x_pow_03 = 16'd178;
        8'd77: x_pow_03 = 16'd179;
        8'd78: x_pow_03 = 16'd179;
        8'd79: x_pow_03 = 16'd180;
        8'd80: x_pow_03 = 16'd181;
        8'd81: x_pow_03 = 16'd181;
        8'd82: x_pow_03 = 16'd182;
        8'd83: x_pow_03 = 16'd183;
        8'd84: x_pow_03 = 16'd183;
        8'd85: x_pow_03 = 16'd184;
        8'd86: x_pow_03 = 16'd185;
        8'd87: x_pow_03 = 16'd185;
        8'd88: x_pow_03 = 16'd186;
        8'd89: x_pow_03 = 16'd187;
        8'd90: x_pow_03 = 16'd187;
        8'd91: x_pow_03 = 16'd188;
        8'd92: x_pow_03 = 16'd189;
        8'd93: x_pow_03 = 16'd189;
        8'd94: x_pow_03 = 16'd190;
        8'd95: x_pow_03 = 16'd190;
        8'd96: x_pow_03 = 16'd191;
        8'd97: x_pow_03 = 16'd192;
        8'd98: x_pow_03 = 16'd192;
        8'd99: x_pow_03 = 16'd193;
        8'd100: x_pow_03 = 16'd193;
        8'd101: x_pow_03 = 16'd194;
        8'd102: x_pow_03 = 16'd194;
        8'd103: x_pow_03 = 16'd195;
        8'd104: x_pow_03 = 16'd196;
        8'd105: x_pow_03 = 16'd196;
        8'd106: x_pow_03 = 16'd197;
        8'd107: x_pow_03 = 16'd197;
        8'd108: x_pow_03 = 16'd198;
        8'd109: x_pow_03 = 16'd198;
        8'd110: x_pow_03 = 16'd199;
        8'd111: x_pow_03 = 16'd199;
        8'd112: x_pow_03 = 16'd200;
        8'd113: x_pow_03 = 16'd201;
        8'd114: x_pow_03 = 16'd201;
        8'd115: x_pow_03 = 16'd202;
        8'd116: x_pow_03 = 16'd202;
        8'd117: x_pow_03 = 16'd203;
        8'd118: x_pow_03 = 16'd203;
        8'd119: x_pow_03 = 16'd204;
        8'd120: x_pow_03 = 16'd204;
        8'd121: x_pow_03 = 16'd205;
        8'd122: x_pow_03 = 16'd205;
        8'd123: x_pow_03 = 16'd206;
        8'd124: x_pow_03 = 16'd206;
        8'd125: x_pow_03 = 16'd207;
        8'd126: x_pow_03 = 16'd207;
        8'd127: x_pow_03 = 16'd208;
        8'd128: x_pow_03 = 16'd208;
        8'd129: x_pow_03 = 16'd209;
        8'd130: x_pow_03 = 16'd209;
        8'd131: x_pow_03 = 16'd210;
        8'd132: x_pow_03 = 16'd210;
        8'd133: x_pow_03 = 16'd211;
        8'd134: x_pow_03 = 16'd211;
        8'd135: x_pow_03 = 16'd212;
        8'd136: x_pow_03 = 16'd212;
        8'd137: x_pow_03 = 16'd212;
        8'd138: x_pow_03 = 16'd213;
        8'd139: x_pow_03 = 16'd213;
        8'd140: x_pow_03 = 16'd214;
        8'd141: x_pow_03 = 16'd214;
        8'd142: x_pow_03 = 16'd215;
        8'd143: x_pow_03 = 16'd215;
        8'd144: x_pow_03 = 16'd216;
        8'd145: x_pow_03 = 16'd216;
        8'd146: x_pow_03 = 16'd217;
        8'd147: x_pow_03 = 16'd217;
        8'd148: x_pow_03 = 16'd217;
        8'd149: x_pow_03 = 16'd218;
        8'd150: x_pow_03 = 16'd218;
        8'd151: x_pow_03 = 16'd219;
        8'd152: x_pow_03 = 16'd219;
        8'd153: x_pow_03 = 16'd220;
        8'd154: x_pow_03 = 16'd220;
        8'd155: x_pow_03 = 16'd220;
        8'd156: x_pow_03 = 16'd221;
        8'd157: x_pow_03 = 16'd221;
        8'd158: x_pow_03 = 16'd222;
        8'd159: x_pow_03 = 16'd222;
        8'd160: x_pow_03 = 16'd223;
        8'd161: x_pow_03 = 16'd223;
        8'd162: x_pow_03 = 16'd223;
        8'd163: x_pow_03 = 16'd224;
        8'd164: x_pow_03 = 16'd224;
        8'd165: x_pow_03 = 16'd225;
        8'd166: x_pow_03 = 16'd225;
        8'd167: x_pow_03 = 16'd225;
        8'd168: x_pow_03 = 16'd226;
        8'd169: x_pow_03 = 16'd226;
        8'd170: x_pow_03 = 16'd227;
        8'd171: x_pow_03 = 16'd227;
        8'd172: x_pow_03 = 16'd227;
        8'd173: x_pow_03 = 16'd228;
        8'd174: x_pow_03 = 16'd228;
        8'd175: x_pow_03 = 16'd229;
        8'd176: x_pow_03 = 16'd229;
        8'd177: x_pow_03 = 16'd229;
        8'd178: x_pow_03 = 16'd230;
        8'd179: x_pow_03 = 16'd230;
        8'd180: x_pow_03 = 16'd231;
        8'd181: x_pow_03 = 16'd231;
        8'd182: x_pow_03 = 16'd231;
        8'd183: x_pow_03 = 16'd232;
        8'd184: x_pow_03 = 16'd232;
        8'd185: x_pow_03 = 16'd233;
        8'd186: x_pow_03 = 16'd233;
        8'd187: x_pow_03 = 16'd233;
        8'd188: x_pow_03 = 16'd234;
        8'd189: x_pow_03 = 16'd234;
        8'd190: x_pow_03 = 16'd234;
        8'd191: x_pow_03 = 16'd235;
        8'd192: x_pow_03 = 16'd235;
        8'd193: x_pow_03 = 16'd235;
        8'd194: x_pow_03 = 16'd236;
        8'd195: x_pow_03 = 16'd236;
        8'd196: x_pow_03 = 16'd237;
        8'd197: x_pow_03 = 16'd237;
        8'd198: x_pow_03 = 16'd237;
        8'd199: x_pow_03 = 16'd238;
        8'd200: x_pow_03 = 16'd238;
        8'd201: x_pow_03 = 16'd238;
        8'd202: x_pow_03 = 16'd239;
        8'd203: x_pow_03 = 16'd239;
        8'd204: x_pow_03 = 16'd239;
        8'd205: x_pow_03 = 16'd240;
        8'd206: x_pow_03 = 16'd240;
        8'd207: x_pow_03 = 16'd240;
        8'd208: x_pow_03 = 16'd241;
        8'd209: x_pow_03 = 16'd241;
        8'd210: x_pow_03 = 16'd242;
        8'd211: x_pow_03 = 16'd242;
        8'd212: x_pow_03 = 16'd242;
        8'd213: x_pow_03 = 16'd243;
        8'd214: x_pow_03 = 16'd243;
        8'd215: x_pow_03 = 16'd243;
        8'd216: x_pow_03 = 16'd244;
        8'd217: x_pow_03 = 16'd244;
        8'd218: x_pow_03 = 16'd244;
        8'd219: x_pow_03 = 16'd245;
        8'd220: x_pow_03 = 16'd245;
        8'd221: x_pow_03 = 16'd245;
        8'd222: x_pow_03 = 16'd246;
        8'd223: x_pow_03 = 16'd246;
        8'd224: x_pow_03 = 16'd246;
        8'd225: x_pow_03 = 16'd247;
        8'd226: x_pow_03 = 16'd247;
        8'd227: x_pow_03 = 16'd247;
        8'd228: x_pow_03 = 16'd248;
        8'd229: x_pow_03 = 16'd248;
        8'd230: x_pow_03 = 16'd248;
        8'd231: x_pow_03 = 16'd249;
        8'd232: x_pow_03 = 16'd249;
        8'd233: x_pow_03 = 16'd249;
        8'd234: x_pow_03 = 16'd249;
        8'd235: x_pow_03 = 16'd250;
        8'd236: x_pow_03 = 16'd250;
        8'd237: x_pow_03 = 16'd250;
        8'd238: x_pow_03 = 16'd251;
        8'd239: x_pow_03 = 16'd251;
        8'd240: x_pow_03 = 16'd251;
        8'd241: x_pow_03 = 16'd252;
        8'd242: x_pow_03 = 16'd252;
        8'd243: x_pow_03 = 16'd252;
        8'd244: x_pow_03 = 16'd253;
        8'd245: x_pow_03 = 16'd253;
        8'd246: x_pow_03 = 16'd253;
        8'd247: x_pow_03 = 16'd254;
        8'd248: x_pow_03 = 16'd254;
        8'd249: x_pow_03 = 16'd254;
        8'd250: x_pow_03 = 16'd254;
        8'd251: x_pow_03 = 16'd255;
        8'd252: x_pow_03 = 16'd255;
        8'd253: x_pow_03 = 16'd255;
        8'd254: x_pow_03 = 16'd256;
        8'd255: x_pow_03 = 16'd256;
        default: x_pow_03 = 16'd0;
    endcase
end

always @(*) begin
    case(y)
        8'd0: y_pow_07 = 16'd0;
        8'd1: y_pow_07 = 16'd5;
        8'd2: y_pow_07 = 16'd9;
        8'd3: y_pow_07 = 16'd11;
        8'd4: y_pow_07 = 16'd14;
        8'd5: y_pow_07 = 16'd16;
        8'd6: y_pow_07 = 16'd19;
        8'd7: y_pow_07 = 16'd21;
        8'd8: y_pow_07 = 16'd23;
        8'd9: y_pow_07 = 16'd25;
        8'd10: y_pow_07 = 16'd27;
        8'd11: y_pow_07 = 16'd28;
        8'd12: y_pow_07 = 16'd30;
        8'd13: y_pow_07 = 16'd32;
        8'd14: y_pow_07 = 16'd34;
        8'd15: y_pow_07 = 16'd35;
        8'd16: y_pow_07 = 16'd37;
        8'd17: y_pow_07 = 16'd38;
        8'd18: y_pow_07 = 16'd40;
        8'd19: y_pow_07 = 16'd42;
        8'd20: y_pow_07 = 16'd43;
        8'd21: y_pow_07 = 16'd45;
        8'd22: y_pow_07 = 16'd46;
        8'd23: y_pow_07 = 16'd48;
        8'd24: y_pow_07 = 16'd49;
        8'd25: y_pow_07 = 16'd50;
        8'd26: y_pow_07 = 16'd52;
        8'd27: y_pow_07 = 16'd53;
        8'd28: y_pow_07 = 16'd55;
        8'd29: y_pow_07 = 16'd56;
        8'd30: y_pow_07 = 16'd57;
        8'd31: y_pow_07 = 16'd59;
        8'd32: y_pow_07 = 16'd60;
        8'd33: y_pow_07 = 16'd61;
        8'd34: y_pow_07 = 16'd62;
        8'd35: y_pow_07 = 16'd64;
        8'd36: y_pow_07 = 16'd65;
        8'd37: y_pow_07 = 16'd66;
        8'd38: y_pow_07 = 16'd68;
        8'd39: y_pow_07 = 16'd69;
        8'd40: y_pow_07 = 16'd70;
        8'd41: y_pow_07 = 16'd71;
        8'd42: y_pow_07 = 16'd72;
        8'd43: y_pow_07 = 16'd74;
        8'd44: y_pow_07 = 16'd75;
        8'd45: y_pow_07 = 16'd76;
        8'd46: y_pow_07 = 16'd77;
        8'd47: y_pow_07 = 16'd78;
        8'd48: y_pow_07 = 16'd80;
        8'd49: y_pow_07 = 16'd81;
        8'd50: y_pow_07 = 16'd82;
        8'd51: y_pow_07 = 16'd83;
        8'd52: y_pow_07 = 16'd84;
        8'd53: y_pow_07 = 16'd85;
        8'd54: y_pow_07 = 16'd86;
        8'd55: y_pow_07 = 16'd87;
        8'd56: y_pow_07 = 16'd89;
        8'd57: y_pow_07 = 16'd90;
        8'd58: y_pow_07 = 16'd91;
        8'd59: y_pow_07 = 16'd92;
        8'd60: y_pow_07 = 16'd93;
        8'd61: y_pow_07 = 16'd94;
        8'd62: y_pow_07 = 16'd95;
        8'd63: y_pow_07 = 16'd96;
        8'd64: y_pow_07 = 16'd97;
        8'd65: y_pow_07 = 16'd98;
        8'd66: y_pow_07 = 16'd99;
        8'd67: y_pow_07 = 16'd100;
        8'd68: y_pow_07 = 16'd101;
        8'd69: y_pow_07 = 16'd103;
        8'd70: y_pow_07 = 16'd104;
        8'd71: y_pow_07 = 16'd105;
        8'd72: y_pow_07 = 16'd106;
        8'd73: y_pow_07 = 16'd107;
        8'd74: y_pow_07 = 16'd108;
        8'd75: y_pow_07 = 16'd109;
        8'd76: y_pow_07 = 16'd110;
        8'd77: y_pow_07 = 16'd111;
        8'd78: y_pow_07 = 16'd112;
        8'd79: y_pow_07 = 16'd113;
        8'd80: y_pow_07 = 16'd114;
        8'd81: y_pow_07 = 16'd115;
        8'd82: y_pow_07 = 16'd116;
        8'd83: y_pow_07 = 16'd117;
        8'd84: y_pow_07 = 16'd118;
        8'd85: y_pow_07 = 16'd119;
        8'd86: y_pow_07 = 16'd120;
        8'd87: y_pow_07 = 16'd121;
        8'd88: y_pow_07 = 16'd122;
        8'd89: y_pow_07 = 16'd123;
        8'd90: y_pow_07 = 16'd123;
        8'd91: y_pow_07 = 16'd124;
        8'd92: y_pow_07 = 16'd125;
        8'd93: y_pow_07 = 16'd126;
        8'd94: y_pow_07 = 16'd127;
        8'd95: y_pow_07 = 16'd128;
        8'd96: y_pow_07 = 16'd129;
        8'd97: y_pow_07 = 16'd130;
        8'd98: y_pow_07 = 16'd131;
        8'd99: y_pow_07 = 16'd132;
        8'd100: y_pow_07 = 16'd133;
        8'd101: y_pow_07 = 16'd134;
        8'd102: y_pow_07 = 16'd135;
        8'd103: y_pow_07 = 16'd136;
        8'd104: y_pow_07 = 16'd137;
        8'd105: y_pow_07 = 16'd138;
        8'd106: y_pow_07 = 16'd138;
        8'd107: y_pow_07 = 16'd139;
        8'd108: y_pow_07 = 16'd140;
        8'd109: y_pow_07 = 16'd141;
        8'd110: y_pow_07 = 16'd142;
        8'd111: y_pow_07 = 16'd143;
        8'd112: y_pow_07 = 16'd144;
        8'd113: y_pow_07 = 16'd145;
        8'd114: y_pow_07 = 16'd146;
        8'd115: y_pow_07 = 16'd147;
        8'd116: y_pow_07 = 16'd147;
        8'd117: y_pow_07 = 16'd148;
        8'd118: y_pow_07 = 16'd149;
        8'd119: y_pow_07 = 16'd150;
        8'd120: y_pow_07 = 16'd151;
        8'd121: y_pow_07 = 16'd152;
        8'd122: y_pow_07 = 16'd153;
        8'd123: y_pow_07 = 16'd154;
        8'd124: y_pow_07 = 16'd155;
        8'd125: y_pow_07 = 16'd155;
        8'd126: y_pow_07 = 16'd156;
        8'd127: y_pow_07 = 16'd157;
        8'd128: y_pow_07 = 16'd158;
        8'd129: y_pow_07 = 16'd159;
        8'd130: y_pow_07 = 16'd160;
        8'd131: y_pow_07 = 16'd161;
        8'd132: y_pow_07 = 16'd161;
        8'd133: y_pow_07 = 16'd162;
        8'd134: y_pow_07 = 16'd163;
        8'd135: y_pow_07 = 16'd164;
        8'd136: y_pow_07 = 16'd165;
        8'd137: y_pow_07 = 16'd166;
        8'd138: y_pow_07 = 16'd167;
        8'd139: y_pow_07 = 16'd167;
        8'd140: y_pow_07 = 16'd168;
        8'd141: y_pow_07 = 16'd169;
        8'd142: y_pow_07 = 16'd170;
        8'd143: y_pow_07 = 16'd171;
        8'd144: y_pow_07 = 16'd172;
        8'd145: y_pow_07 = 16'd172;
        8'd146: y_pow_07 = 16'd173;
        8'd147: y_pow_07 = 16'd174;
        8'd148: y_pow_07 = 16'd175;
        8'd149: y_pow_07 = 16'd176;
        8'd150: y_pow_07 = 16'd177;
        8'd151: y_pow_07 = 16'd177;
        8'd152: y_pow_07 = 16'd178;
        8'd153: y_pow_07 = 16'd179;
        8'd154: y_pow_07 = 16'd180;
        8'd155: y_pow_07 = 16'd181;
        8'd156: y_pow_07 = 16'd181;
        8'd157: y_pow_07 = 16'd182;
        8'd158: y_pow_07 = 16'd183;
        8'd159: y_pow_07 = 16'd184;
        8'd160: y_pow_07 = 16'd185;
        8'd161: y_pow_07 = 16'd186;
        8'd162: y_pow_07 = 16'd186;
        8'd163: y_pow_07 = 16'd187;
        8'd164: y_pow_07 = 16'd188;
        8'd165: y_pow_07 = 16'd189;
        8'd166: y_pow_07 = 16'd190;
        8'd167: y_pow_07 = 16'd190;
        8'd168: y_pow_07 = 16'd191;
        8'd169: y_pow_07 = 16'd192;
        8'd170: y_pow_07 = 16'd193;
        8'd171: y_pow_07 = 16'd194;
        8'd172: y_pow_07 = 16'd194;
        8'd173: y_pow_07 = 16'd195;
        8'd174: y_pow_07 = 16'd196;
        8'd175: y_pow_07 = 16'd197;
        8'd176: y_pow_07 = 16'd197;
        8'd177: y_pow_07 = 16'd198;
        8'd178: y_pow_07 = 16'd199;
        8'd179: y_pow_07 = 16'd200;
        8'd180: y_pow_07 = 16'd201;
        8'd181: y_pow_07 = 16'd201;
        8'd182: y_pow_07 = 16'd202;
        8'd183: y_pow_07 = 16'd203;
        8'd184: y_pow_07 = 16'd204;
        8'd185: y_pow_07 = 16'd204;
        8'd186: y_pow_07 = 16'd205;
        8'd187: y_pow_07 = 16'd206;
        8'd188: y_pow_07 = 16'd207;
        8'd189: y_pow_07 = 16'd208;
        8'd190: y_pow_07 = 16'd208;
        8'd191: y_pow_07 = 16'd209;
        8'd192: y_pow_07 = 16'd210;
        8'd193: y_pow_07 = 16'd211;
        8'd194: y_pow_07 = 16'd211;
        8'd195: y_pow_07 = 16'd212;
        8'd196: y_pow_07 = 16'd213;
        8'd197: y_pow_07 = 16'd214;
        8'd198: y_pow_07 = 16'd214;
        8'd199: y_pow_07 = 16'd215;
        8'd200: y_pow_07 = 16'd216;
        8'd201: y_pow_07 = 16'd217;
        8'd202: y_pow_07 = 16'd217;
        8'd203: y_pow_07 = 16'd218;
        8'd204: y_pow_07 = 16'd219;
        8'd205: y_pow_07 = 16'd220;
        8'd206: y_pow_07 = 16'd220;
        8'd207: y_pow_07 = 16'd221;
        8'd208: y_pow_07 = 16'd222;
        8'd209: y_pow_07 = 16'd223;
        8'd210: y_pow_07 = 16'd223;
        8'd211: y_pow_07 = 16'd224;
        8'd212: y_pow_07 = 16'd225;
        8'd213: y_pow_07 = 16'd226;
        8'd214: y_pow_07 = 16'd226;
        8'd215: y_pow_07 = 16'd227;
        8'd216: y_pow_07 = 16'd228;
        8'd217: y_pow_07 = 16'd229;
        8'd218: y_pow_07 = 16'd229;
        8'd219: y_pow_07 = 16'd230;
        8'd220: y_pow_07 = 16'd231;
        8'd221: y_pow_07 = 16'd232;
        8'd222: y_pow_07 = 16'd232;
        8'd223: y_pow_07 = 16'd233;
        8'd224: y_pow_07 = 16'd234;
        8'd225: y_pow_07 = 16'd235;
        8'd226: y_pow_07 = 16'd235;
        8'd227: y_pow_07 = 16'd236;
        8'd228: y_pow_07 = 16'd237;
        8'd229: y_pow_07 = 16'd237;
        8'd230: y_pow_07 = 16'd238;
        8'd231: y_pow_07 = 16'd239;
        8'd232: y_pow_07 = 16'd240;
        8'd233: y_pow_07 = 16'd240;
        8'd234: y_pow_07 = 16'd241;
        8'd235: y_pow_07 = 16'd242;
        8'd236: y_pow_07 = 16'd242;
        8'd237: y_pow_07 = 16'd243;
        8'd238: y_pow_07 = 16'd244;
        8'd239: y_pow_07 = 16'd245;
        8'd240: y_pow_07 = 16'd245;
        8'd241: y_pow_07 = 16'd246;
        8'd242: y_pow_07 = 16'd247;
        8'd243: y_pow_07 = 16'd248;
        8'd244: y_pow_07 = 16'd248;
        8'd245: y_pow_07 = 16'd249;
        8'd246: y_pow_07 = 16'd250;
        8'd247: y_pow_07 = 16'd250;
        8'd248: y_pow_07 = 16'd251;
        8'd249: y_pow_07 = 16'd252;
        8'd250: y_pow_07 = 16'd252;
        8'd251: y_pow_07 = 16'd253;
        8'd252: y_pow_07 = 16'd254;
        8'd253: y_pow_07 = 16'd255;
        8'd254: y_pow_07 = 16'd255;
        8'd255: y_pow_07 = 16'd256;
        default: y_pow_07 = 16'd0;
    endcase
end
endmodule
